module top_module( 
    input a,b,c,
    output w,x,y,z );

endmodule